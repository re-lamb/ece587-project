/*
 * ECE587 Fall 2024 Final Project
 * R.E. Lamb
 *
 * CPU top level 
 */
`include "defs.svh"

module sim(
  );
  
  /*
  memory mem(         - 95%
  );
  
  fetch ifu(          - 95%
  );
  
  bpred bp(           - 0% - xxx
  );
  
  decode id(          - 75% - needs rob_packet/fu_select
  );
  
  reorder rob(        - 0%
  );
  
  freelist fl(        - 85% - needs freelist_t/rollback
  );
  
  maptable rmap(      - 85% - copy mem/regfile, needs rollback
  );
  
  regfile regs(       - 95%
  );
  
  issue is(           - 0% - use logisim design
  );
  
  loadstore lsu(      - 0% - xxx
  );
  
  alu alu(            - 0% - recycle
  );
  
  branch bru(         - 0% - simple
  );
  */
  
endmodule
